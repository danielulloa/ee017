* Con est� sintaxis LTspice pone
* autom�ticamente el par�metro per�odo
* En el s�mbolo y queda funcionando perfectamente.
* Luego se reacomoda el dibujo seg�n nuestras necesidades
*
.subckt promediador ent sal
+periodo=1ms
T1 ent 0 vdemorada 0 Td={periodo} Z0=1g
R1 vdemorada 0 1g
G1 0 sal ent vdemorada 1
C1 sal 0 {periodo} ic=0 Rser=0 Lser=0 Rpar=1g Cpar=0
.ends promediador
