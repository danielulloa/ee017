* LF411C OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* http://www.ti.com/product/LF411
* CREATED USING PARTS RELEASE 4.01 ON 06/27/89 AT 08:19
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT LF411C   1 2 3 4 5
*
  C1   11 12 3.498E-12
  C2    6  7 15.00E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  FB    7 99 POLY(5) VB VC VE VLP VLN 0 28.29E6 -30E6 30E6 30E6 -30E6
  GA    6  0 11 12 282.8E-6
  GCM   0  6 10 99 1.590E-9
  ISS   3 10 DC 195.0E-6
  HLIM 90  0 VLIM 1K
  J1   11  2 10 JX
  J2   12  1 10 JX
  R2    6  9 100.0E3
  RD1   4 11 3.536E3
  RD2   4 12 3.536E3
  RO1   8  5 50
  RO2   7 99 25
  RP    3  4 15.00E3
  RSS  10 99 1.026E6
  VB    9  0 DC 0
  VC    3 53 DC 2.200
  VE   54  4 DC 2.200
  VLIM  7  8 DC 0
  VLP  91  0 DC 30
  VLN   0 92 DC 30
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=12.50E-12 BETA=250.1E-6 VTO=-1)
.ENDS
